module top(input A, input B, output SUM);
  assign SUM = A ^ B;  // Simple XOR gate
endmodule
